****AND_Gate circuit design****
