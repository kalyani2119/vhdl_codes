# vhdl_codes
  ****NOT_GATE circuit design****
  
